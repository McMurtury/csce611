module CSCE611_regfile_testbench(

input CLOCK_50,

output [3:0] tiamat
);

endmodule
